library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_led is

  port (
	INIT_DONE : out std_logic;
	LVDS23n : out std_logic;
	LVDS22p : out std_logic;
	LVDS22n : out std_logic;
	VREF0B1 : out std_logic;
	PIN_6 : out std_logic;
	LVDS21p : out std_logic;
	LVDS21n : out std_logic;
	DPCLK1 : out std_logic;
	LVDS20p : out std_logic;
	LVDS20n : out std_logic;
	LVDS19p : out std_logic;
	LVDS19n : out std_logic;
	LVDS18p : out std_logic;
	LVDS18n : out std_logic;
	LVDS17p : out std_logic;
	LVDS17n : out std_logic;
	LVDS16p : out std_logic;
	LVDS16n : out std_logic;
	VREF1B1 : out std_logic;
	nCSO : out std_logic;
	CLK0 : in std_logic;
	CLK1 : in std_logic;
	ASDO : out std_logic;
	PLL1_OUTp : out std_logic;
	PLL1_OUTn : out std_logic;
	LVDS7n : out std_logic;
	LVDS6p : out std_logic;
	LVDS6n : out std_logic;
	LVDS5p : out std_logic;
	LVDS5n : out std_logic;
	LVDS4p : out std_logic;
	LVDS4n : out std_logic;
	LVDS3p : out std_logic;
	LVDS3n : out std_logic;
	DPCLK0 : out std_logic;
	LVDS2p : out std_logic;
	LVDS2n : out std_logic;
	PIN_56 : out std_logic;
	LVDS1p : out std_logic;
	LVDS1n : out std_logic;
	LVDS0p : out std_logic;
	LVDS0n : out std_logic;
	LVDS102p : out std_logic;
	LVDS102n : out std_logic;
	LVDS101p : out std_logic;
	LVDS101n : out std_logic;
	LVDS100p : out std_logic;
	LVDS100n : out std_logic;
	LVDS99p  : out std_logic;
	LVDS99n  : out std_logic;
	DPCLK7   : out std_logic;
	LVDS98p  : out std_logic;
	LVDS98n  : out std_logic;
	LVDS97p  : out std_logic;
	LVDS97n  : out std_logic;
	LVDS96p  : out std_logic;
	LVDS95p  : out std_logic;
	LVDS95n  : out std_logic;
	LVDS94p  : out std_logic;
	LVDS94n  : out std_logic;
	LVDS93p  : out std_logic;
	LVDS93n  : out std_logic;
	LVDS92p  : out std_logic;
	LVDS87p  : out std_logic;
	LVDS87n  : out std_logic;
	LVDS86p  : out std_logic;
	LVDS86n  : out std_logic;
	LVDS85p  : out std_logic;
	LVDS85n  : out std_logic;
	LVDS80p  : out std_logic;
	LVDS80n  : out std_logic;
	PIN_106  : out std_logic;
	DPCLK6   : out std_logic;
	LVDS79p  : out std_logic;
	LVDS79n  : out std_logic;
	LVDS78p  : out std_logic;
	LVDS78n  : out std_logic;
	LVDS77p  : out std_logic;
	LVDS77n  : out std_logic;
	LVDS76p  : out std_logic;
	LVDS76n  : out std_logic;
	LVDS75n  : out std_logic;
	LVDS75p  : out std_logic;
	LVDS74n  : out std_logic;
	LVDS74p  : out std_logic;
	LVDS73n  : out std_logic;
	LVDS73p  : out std_logic;
	PIN_128  : out std_logic;
	DPCLK5   : out std_logic;
	LVDS72n  : out std_logic;
	LVDS72p  : out std_logic;
	LVDS71n  : out std_logic;
	LVDS71p  : out std_logic;
	LVDS70n  : out std_logic;
	LVDS70p  : out std_logic;
	LVDS69n  : out std_logic;
	LVDS69p  : out std_logic;
	LVDS68n  : out std_logic;
	LVDS68p  : out std_logic;
	PLL2_OUTn : out std_logic;
	PLL2_OUTp : out std_logic;
	CLK3  : in std_logic;
	CLK2  : in std_logic;
	LVDS59n  : out std_logic;
	LVDS59p  : out std_logic;
	LVDS58n  : out std_logic;
	LVDS58p  : out std_logic;
	LVDS57n  : out std_logic;
	LVDS57p  : out std_logic;
	LVDS56n  : out std_logic;
	LVDS56p  : out std_logic;
	LVDS55n  : out std_logic;
	LVDS55p  : out std_logic;
	LVDS54n  : out std_logic;
	LVDS54p  : out std_logic;
	DPCLK4  : out std_logic;
	LVDS53n  : out std_logic;
	LVDS53p  : out std_logic;
	PIN_175  : out std_logic;
	LVDS52n  : out std_logic;
	LVDS52p  : out std_logic;
	LVDS51n  : out std_logic;
	LVDS51p  : out std_logic;
	LVDS50n  : out std_logic;
	LVDS50p  : out std_logic;
	LVDS49n  : out std_logic;
	LVDS49p  : out std_logic;
	LVDS48n  : out std_logic;
	LVDS48p  : out std_logic;
	LVDS47n  : out std_logic;
	LVDS47p  : out std_logic;
	DPCLK3  : out std_logic;
	PIN_195  : out std_logic;
	LVDS46n  : out std_logic;
	LVDS46p  : out std_logic;
	LVDS41n  : out std_logic;
	LVDS41p  : out std_logic;
	LVDS40n  : out std_logic;
	LVDS40p  : out std_logic;
	LVDS39n  : out std_logic;
	LVDS39p  : out std_logic;
	LVDS34p  : out std_logic;
	LVDS33n  : out std_logic;
	LVDS33p  : out std_logic;
	LVDS32n  : out std_logic;
	LVDS32p  : out std_logic;
	LVDS31n  : out std_logic;
	LVDS31p  : out std_logic;
	LVDS30p  : out std_logic;
	LVDS29n  : out std_logic;
	LVDS29p  : out std_logic;
	LVDS28n  : out std_logic;
	LVDS28p  : out std_logic;
	DPCLK2  : out std_logic;
	LVDS27n  : out std_logic;
	LVDS27p  : out std_logic;
	LVDS26n  : out std_logic;
	LVDS26p  : out std_logic;
	LVDS25n  : out std_logic;
	LVDS25p  : out std_logic;
	LVDS24n  : out std_logic;
	LVDS24p  : out std_logic
    );

end test_led;

architecture behaviour of test_led is
begin
	INIT_DONE <= '1';
	LVDS23n <= '1';
	LVDS22p <= '1';
	LVDS22n <= '1';
	VREF0B1 <= '1';
	PIN_6 <= '1';
	LVDS21p <= '1';
	LVDS21n <= '1';
	DPCLK1 <= '1';
	LVDS20p <= '1';
	LVDS20n <= '1';
	LVDS19p <= '1';
	LVDS19n <= '1';
	LVDS18p <= '1';
	LVDS18n <= '1';
	LVDS17p <= '1';
	LVDS17n <= '1';
	LVDS16p <= '1';
	LVDS16n <= '1';
	VREF1B1 <= '1';
	nCSO <= '1';
	ASDO <= '1';
	PLL1_OUTp <= '1';
	PLL1_OUTn <= '1';
	LVDS7n <= '1';
	LVDS6p <= '1';
	LVDS6n <= '1';
	LVDS5p <= '1';
	LVDS5n <= '1';
	LVDS4p <= '1';
	LVDS4n <= '1';
	LVDS3p <= '1';
	LVDS3n <= '1';
	DPCLK0 <= '1';
	LVDS2p <= '1';
	LVDS2n <= '1';
	PIN_56 <= '1';
	LVDS1p <= '1';
	LVDS1n <= '1';
	LVDS0p <= '1';
	LVDS0n <= '1';
	LVDS102p <= '1';
	LVDS102n <= '1';
	LVDS101p <= '1';
	LVDS101n <= '1';
	LVDS100p <= '1';
	LVDS100n <= '1';
	LVDS99p  <= '1';
	LVDS99n  <= '1';
	DPCLK7   <= '1';
	LVDS98p  <= '1';
	LVDS98n  <= '1';
	LVDS97p  <= '1';
	LVDS97n  <= '1';
	LVDS96p  <= '1';
	LVDS95p  <= '1';
	LVDS95n  <= '1';
	LVDS94p  <= '1';
	LVDS94n  <= '1';
	LVDS93p  <= '1';
	LVDS93n  <= '1';
	LVDS92p  <= '1';
	LVDS87p  <= '1';
	LVDS87n  <= '1';
	LVDS86p  <= '1';
	LVDS86n  <= '1';
	LVDS85p  <= '1';
	LVDS85n  <= '1';
	LVDS80p  <= '1';
	LVDS80n  <= '1';
	PIN_106  <= '1';
	DPCLK6   <= '1';
	LVDS79p  <= '1';
	LVDS79n  <= '1';
	LVDS78p  <= '1';
	LVDS78n  <= '1';
	LVDS77p  <= '1';
	LVDS77n  <= '1';
	LVDS76p  <= '1';
	LVDS76n  <= '1';
	LVDS75n  <= '1';
	LVDS75p  <= '1';
	LVDS74n  <= '1';
	LVDS74p  <= '1';
	LVDS73n  <= '1';
	LVDS73p  <= '1';
	PIN_128  <= '1';
	DPCLK5   <= '1';
	LVDS72n  <= '1';
	LVDS72p  <= '1';
	LVDS71n  <= '1';
	LVDS71p  <= '1';
	LVDS70n  <= '1';
	LVDS70p  <= '1';
	LVDS69n  <= '1';
	LVDS69p  <= '1';
	LVDS68n  <= '1';
	LVDS68p  <= '1';
	PLL2_OUTn <= '1';
	PLL2_OUTp <= '1';
	LVDS59n  <= '1';
	LVDS59p  <= '1';
	LVDS58n  <= '1';
	LVDS58p  <= '1';
	LVDS57n  <= '1';
	LVDS57p  <= '1';
	LVDS56n  <= '1';
	LVDS56p  <= '1';
	LVDS55n  <= '1';
	LVDS55p  <= '1';
	LVDS54n  <= '1';
	LVDS54p  <= '1';
	DPCLK4  <= '1';
	LVDS53n  <= '1';
	LVDS53p  <= '1';
	PIN_175  <= '1';
	LVDS52n  <= '1';
	LVDS52p  <= '1';
	LVDS51n  <= '1';
	LVDS51p  <= '1';
	LVDS50n  <= '1';
	LVDS50p  <= '1';
	LVDS49n  <= '1';
	LVDS49p  <= '1';
	LVDS48n  <= '1';
	LVDS48p  <= '1';
	LVDS47n  <= '1';
	LVDS47p  <= '1';
	DPCLK3  <= '1';
	PIN_195  <= '1';
	LVDS46n  <= '1';
	LVDS46p  <= '1';
	LVDS41n  <= '1';
	LVDS41p  <= '1';
	LVDS40n  <= '1';
	LVDS40p  <= '1';
	LVDS39n  <= '1';
	LVDS39p  <= '1';
	LVDS34p  <= '1';
	LVDS33n  <= '1';
	LVDS33p  <= '1';
	LVDS32n  <= '1';
	LVDS32p  <= '1';
	LVDS31n  <= '1';
	LVDS31p  <= '1';
	LVDS30p  <= '1';
	LVDS29n  <= '1';
	LVDS29p  <= '1';
	LVDS28n  <= '1';
	LVDS28p  <= '1';
	DPCLK2  <= '1';
	LVDS27n  <= '1';
	LVDS27p  <= '1';
	LVDS26n  <= '1';
	LVDS26p  <= '1';
	LVDS25n  <= '1';
	LVDS25p  <= '1';
	LVDS24n  <= '1';
	LVDS24p  <= '1';	
end behaviour;